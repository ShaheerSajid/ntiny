`define PWM_PRESCALER_REG 8'h00
`define PWM_CONTROL_REG   8'h01 
`define PWM_PERIOD1_REG    8'h02
`define PWM_PERIOD2_REG    8'h03 
`define PWM_COMPARE1_REG   8'h04
`define PWM_COMPARE2_REG   8'h05 
`define PWM_DEADTIME1_REG   8'h06 
`define PWM_DEADTIME2_REG   8'h07 




