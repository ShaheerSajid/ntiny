`define PRESCALAR_REG 32'h00
`define COUNT_REG     32'h01
`define CONTROL_REG   32'h02
`define STATUS_REG    32'h03
`define COMPARE_REG   32'h04