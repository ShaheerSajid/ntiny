module zba_zbb (
	
	input[31:0] in1_i,
				in2_i, 
	output logic[31:0]  out_sh1_add_o,
						out_sh2_add_o,
						out_sh3_add_o,
						out_clz_o,
						out_ctz_o,
						out_andn_o,
						out_orn_o,
						out_xnor_o,
						out_orc_o,
						out_rev8_o,
						out_cpop_o,
						out_min_o,
						out_max_o,
						out_minu_o,
						out_maxu_o,
						out_sextb_o,
						out_sexth_o,
						out_zexth_o,
						out_rol_o,
						out_ror_o
				);


integer i;
wire logic temp_cond; 
wire logic temp_cond_s; 

always_comb
	begin
		casez (in1_i)
				32'b00000000000000000000000000000000: out_clz_o = 32'd32;
				32'b00000000000000000000000000000001: out_clz_o = 32'd31;
				32'b0000000000000000000000000000001?: out_clz_o = 32'd30;
				32'b000000000000000000000000000001??: out_clz_o = 32'd29;
				32'b00000000000000000000000000001???: out_clz_o = 32'd28;
				32'b0000000000000000000000000001????: out_clz_o = 32'd27;
				32'b000000000000000000000000001?????: out_clz_o = 32'd26;
				32'b00000000000000000000000001??????: out_clz_o = 32'd25;
				32'b0000000000000000000000001???????: out_clz_o = 32'd24;
				32'b000000000000000000000001????????: out_clz_o = 32'd23;
				32'b00000000000000000000001?????????: out_clz_o = 32'd22;
				32'b0000000000000000000001??????????: out_clz_o = 32'd21;
				32'b000000000000000000001???????????: out_clz_o = 32'd20;
				32'b00000000000000000001????????????: out_clz_o = 32'd19;
				32'b0000000000000000001?????????????: out_clz_o = 32'd18;
				32'b000000000000000001??????????????: out_clz_o = 32'd17;
				32'b00000000000000001???????????????: out_clz_o = 32'd16;
				32'b0000000000000001????????????????: out_clz_o = 32'd15;
				32'b000000000000001?????????????????: out_clz_o = 32'd14;
				32'b00000000000001??????????????????: out_clz_o = 32'd13;
				32'b0000000000001???????????????????: out_clz_o = 32'd12;
				32'b000000000001????????????????????: out_clz_o = 32'd11;
				32'b00000000001?????????????????????: out_clz_o = 32'd10;
				32'b0000000001??????????????????????: out_clz_o = 32'd9;
				32'b000000001???????????????????????: out_clz_o = 32'd8;
				32'b00000001????????????????????????: out_clz_o = 32'd7;
				32'b0000001?????????????????????????: out_clz_o = 32'd6;
				32'b000001??????????????????????????: out_clz_o = 32'd5;
				32'b00001???????????????????????????: out_clz_o = 32'd4;
				32'b0001????????????????????????????: out_clz_o = 32'd3;
				32'b001?????????????????????????????: out_clz_o = 32'd2;
				32'b01??????????????????????????????: out_clz_o = 32'd1;
				32'b1???????????????????????????????: out_clz_o = 32'd0;
				default: out_clz_o = 32'd0;
		endcase
		
		casez (in1_i)
				32'b???????????????????????????????1: out_ctz_o = 32'd0;
				32'b??????????????????????????????10: out_ctz_o = 32'd1;
				32'b?????????????????????????????100: out_ctz_o = 32'd2;
				32'b????????????????????????????1000: out_ctz_o = 32'd3;
				32'b???????????????????????????10000: out_ctz_o = 32'd4;
				32'b??????????????????????????100000: out_ctz_o = 32'd5;
				32'b?????????????????????????1000000: out_ctz_o = 32'd6;
				32'b????????????????????????10000000: out_ctz_o = 32'd7;
				32'b???????????????????????100000000: out_ctz_o = 32'd8;
				32'b??????????????????????1000000000: out_ctz_o = 32'd9;
				32'b?????????????????????10000000000: out_ctz_o = 32'd10;
				32'b????????????????????100000000000: out_ctz_o = 32'd11;
				32'b???????????????????1000000000000: out_ctz_o = 32'd12;
				32'b??????????????????10000000000000: out_ctz_o = 32'd13;
				32'b?????????????????100000000000000: out_ctz_o = 32'd14;
				32'b????????????????1000000000000000: out_ctz_o = 32'd15;
				32'b???????????????10000000000000000: out_ctz_o = 32'd16;
				32'b??????????????100000000000000000: out_ctz_o = 32'd17;
				32'b?????????????1000000000000000000: out_ctz_o = 32'd18;
				32'b????????????10000000000000000000: out_ctz_o = 32'd19;
				32'b???????????100000000000000000000: out_ctz_o = 32'd20;
				32'b??????????1000000000000000000000: out_ctz_o = 32'd21;
				32'b?????????10000000000000000000000: out_ctz_o = 32'd22;
				32'b????????100000000000000000000000: out_ctz_o = 32'd23;
				32'b???????1000000000000000000000000: out_ctz_o = 32'd24;
				32'b??????10000000000000000000000000: out_ctz_o = 32'd25;
				32'b?????100000000000000000000000000: out_ctz_o = 32'd26;
				32'b????1000000000000000000000000000: out_ctz_o = 32'd27;
				32'b???10000000000000000000000000000: out_ctz_o = 32'd28;
				32'b??100000000000000000000000000000: out_ctz_o = 32'd29;
				32'b?1000000000000000000000000000000: out_ctz_o = 32'd30;
				32'b10000000000000000000000000000000: out_ctz_o = 32'd31;
				32'b00000000000000000000000000000000: out_ctz_o = 32'd32;
				default: out_ctz_o = 32'd0;
		endcase
end
/****************************************adder tree *********************/
var logic[2:0] stage1 [15:0];
var logic[3:0] stage2 [7:0];
var logic[4:0] stage3 [3:0];
var logic[5:0] stage4 [1:0];

always_comb
begin
	out_cpop_o =0;
	for (i =0 ;i<16 ;i= i+1 ) begin		//adder tree first stage
		stage1[i] = in1_i[2*i] + in1_i[2*i + 1]; 	
	end

	for (i =0 ;i<8 ;i= i+1 ) begin		//adder tree second stage
		stage2[i] = stage1[2*i] + stage1[2*i + 1]; 	
	end
	
	for (i =0 ;i<4 ;i= i+1 ) begin		//adder tree third stage
		stage3[i] = stage2[2*i] + stage2[2*i + 1]; 	
	end

	for (i =0 ;i<2 ;i= i+1 ) begin		//adder tree fourth stage
		stage4[i] = stage3[2*i] + stage3[2*i + 1]; 	
	end
	out_cpop_o = stage4[0] + stage4[1];
end

/************shift and add*****************************************/
assign out_sh1_add_o = in2_i + (in1_i << 1);
assign out_sh2_add_o = in2_i + (in1_i << 2);
assign out_sh3_add_o = in2_i + (in1_i << 3);
/************ Logical with Not ************************************/ 
always_comb
begin
out_andn_o = in1_i&~in2_i;
out_orn_o = in1_i|~in2_i;
out_xnor_o = ~(in1_i^in2_i);
end
/****************** Min/max Instructions ********************/
assign temp_cond = in1_i < in2_i;
assign out_minu_o = temp_cond? in1_i:in2_i;
assign out_maxu_o = temp_cond? in2_i:in1_i;

assign temp_cond_s = $signed(in1_i) < $signed(in2_i);
assign out_min_o = temp_cond_s? in1_i:in2_i;
assign out_max_o = temp_cond_s? in2_i:in1_i;
/******** Sign Extend ***************/
assign out_sextb_o = {{24{in1_i[7]}},in1_i[7:0]};
assign out_sexth_o = {{16{in1_i[15]}},in1_i[15:0]};
assign out_zexth_o = {16'd0,in1_i[15:0]};
/******************* Bitwise rotation ************************/
assign out_ror_o = (in1_i >> in2_i[4:0]) | (in1_i << (32 - in2_i[4:0]));
assign out_rol_o = (in1_i << in2_i[4:0]) | (in1_i >> (32 - in2_i[4:0]));
/************** out_orc_o **************/
always_comb
begin
	out_orc_o[7:0] = {8{|(in1_i[7:0])}};
	out_orc_o[15:8] = {8{|(in1_i[15:8])}};
	out_orc_o[23:16] = {8{|(in1_i[23:16])}};
	out_orc_o[31:24] = {8{|(in1_i[31:24])}};
end
/******************************** Byte-reverse *********************/
always_comb
begin
	out_rev8_o[7:0] = in1_i[31:24];
	out_rev8_o[15:8] = in1_i[23:16];
	out_rev8_o[23:16] = in1_i[15:8];
	out_rev8_o[31:24] = in1_i[7:0];
end

endmodule 



